module InstructMem(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	case(Address[30:2])	//Address Must Be Word Aligned.
		0: Instruction <= 32'b00001000000000000000000000000011;
		1: Instruction <= 32'b00001000000000000000000001010011;
		2: Instruction <= 32'b00001000000000000000000001111100;
		3: Instruction <= 32'b00111100000100010100000000000000;
		4: Instruction <= 32'b00111100000111010000000000000000;
		5: Instruction <= 32'b00100011101111010000001111111100;
		6: Instruction <= 32'b00111100000100100000000000000000;
		7: Instruction <= 32'b00100000000010010000000001000000;
		8: Instruction <= 32'b10101110010010010000000000000000;
		9: Instruction <= 32'b00100000000010010000000001111001;
		10: Instruction <= 32'b10101110010010010000000000000100;
		11: Instruction <= 32'b00100000000010010000000000100100;
		12: Instruction <= 32'b10101110010010010000000000001000;
		13: Instruction <= 32'b00100000000010010000000000110000;
		14: Instruction <= 32'b10101110010010010000000000001100;
		15: Instruction <= 32'b00100000000010010000000000011001;
		16: Instruction <= 32'b10101110010010010000000000010000;
		17: Instruction <= 32'b00100000000010010000000000010010;
		18: Instruction <= 32'b10101110010010010000000000010100;
		19: Instruction <= 32'b00100000000010010000000000000010;
		20: Instruction <= 32'b10101110010010010000000000011000;
		21: Instruction <= 32'b00100000000010010000000001111000;
		22: Instruction <= 32'b10101110010010010000000000011100;
		23: Instruction <= 32'b00100000000010010000000000000000;
		24: Instruction <= 32'b10101110010010010000000000100000;
		25: Instruction <= 32'b00100000000010010000000000010000;
		26: Instruction <= 32'b10101110010010010000000000100100;
		27: Instruction <= 32'b00100000000010010000000000001000;
		28: Instruction <= 32'b10101110010010010000000000101000;
		29: Instruction <= 32'b00100000000010010000000000000011;
		30: Instruction <= 32'b10101110010010010000000000101100;
		31: Instruction <= 32'b00100000000010010000000001000110;
		32: Instruction <= 32'b10101110010010010000000000110000;
		33: Instruction <= 32'b00100000000010010000000000100001;
		34: Instruction <= 32'b10101110010010010000000000110100;
		35: Instruction <= 32'b00100000000010010000000000000110;
		36: Instruction <= 32'b10101110010010010000000000111000;
		37: Instruction <= 32'b00100000000010010000000000001110;
		38: Instruction <= 32'b10101110010010010000000000111100;
		39: Instruction <= 32'b00111100000010010000000000000000;
		40: Instruction <= 32'b10101110001010010000000000001000;
		41: Instruction <= 32'b00111100000010100000000000000000;
		42: Instruction <= 32'b00100001001010101111111110000000;
		43: Instruction <= 32'b10101110001010100000000000000000;
		44: Instruction <= 32'b00111100000010010000000000000000;
		45: Instruction <= 32'b00100001001010011111111100000000;
		46: Instruction <= 32'b10101110001010010000000000000100;
		47: Instruction <= 32'b00111100000010010000000000000000;
		48: Instruction <= 32'b00100001001010010000000000000011;
		49: Instruction <= 32'b10101110001010010000000000001000;
		50: Instruction <= 32'b00111100000010100000000000000000;
		51: Instruction <= 32'b00100001010010100000000000010011;
		52: Instruction <= 32'b10101110001010100000000000100000;
		53: Instruction <= 32'b10001110001010100000000000100000;
		54: Instruction <= 32'b00110001010010010000000000001000;
		55: Instruction <= 32'b00010001001000001111111111111101;
		56: Instruction <= 32'b10001110001101010000000000011100;
		57: Instruction <= 32'b10001110001010100000000000100000;
		58: Instruction <= 32'b00110001010010010000000000001000;
		59: Instruction <= 32'b00010001001000001111111111111101;
		60: Instruction <= 32'b10001110001101100000000000011100;
		61: Instruction <= 32'b00000000000101010010000000100000;
		62: Instruction <= 32'b00000000000101100010100000100000;
		63: Instruction <= 32'b00001100000000000000000001000011;
		64: Instruction <= 32'b10101110001000100000000000011000;
		65: Instruction <= 32'b10101110001000100000000000001100;
		66: Instruction <= 32'b00001000000000000000000001000010;
		67: Instruction <= 32'b00000000100001010100100000101010;
		68: Instruction <= 32'b00010001001000000000000000000011;
		69: Instruction <= 32'b00000000000001010101000000100000;
		70: Instruction <= 32'b00000000000001000010100000100000;
		71: Instruction <= 32'b00000000000010100010000000100000;
		72: Instruction <= 32'b00010000101000000000000000001000;
		73: Instruction <= 32'b00000000100001010100100000101010;
		74: Instruction <= 32'b00010101001000000000000000000010;
		75: Instruction <= 32'b00000000100001010010000000100010;
		76: Instruction <= 32'b00001000000000000000000001001001;
		77: Instruction <= 32'b00000000000001010101000000100000;
		78: Instruction <= 32'b00000000000001000010100000100000;
		79: Instruction <= 32'b00000000000010100010000000100000;
		80: Instruction <= 32'b00001000000000000000000001001000;
		81: Instruction <= 32'b00000000000001000001000000100000;
		82: Instruction <= 32'b00000011111000000000000000001000;
		83: Instruction <= 32'b00100011101111011111111111110100;
		84: Instruction <= 32'b10101111101010010000000000000000;
		85: Instruction <= 32'b10101111101010100000000000000100;
		86: Instruction <= 32'b10101111101010110000000000001000;
		87: Instruction <= 32'b00111100000010010000000000000000;
		88: Instruction <= 32'b00100001001010010000000000000001;
		89: Instruction <= 32'b10101110001010010000000000001000;
		90: Instruction <= 32'b00110010101010010000000000001111;
		91: Instruction <= 32'b00000000000010010100100010000000;
		92: Instruction <= 32'b00000001001100100101000000100000;
		93: Instruction <= 32'b10001101010010110000000000000000;
		94: Instruction <= 32'b00100001011010110000000100000000;
		95: Instruction <= 32'b10101110001010110000000000010100;
		96: Instruction <= 32'b00110010101010010000000011110000;
		97: Instruction <= 32'b00000000000010010100100010000010;
		98: Instruction <= 32'b00000001001100100101000000100000;
		99: Instruction <= 32'b10001101010010110000000000000000;
		100: Instruction <= 32'b00100001011010110000001000000000;
		101: Instruction <= 32'b10101110001010110000000000010100;
		102: Instruction <= 32'b00110010110010010000000000001111;
		103: Instruction <= 32'b00000000000010010100100010000000;
		104: Instruction <= 32'b00000001001100100101000000100000;
		105: Instruction <= 32'b10001101010010110000000000000000;
		106: Instruction <= 32'b00100001011010110000010000000000;
		107: Instruction <= 32'b10101110001010110000000000010100;
		108: Instruction <= 32'b00110010110010010000000011110000;
		109: Instruction <= 32'b00000000000010010100100010000010;
		110: Instruction <= 32'b00000001001100100101000000100000;
		111: Instruction <= 32'b10001101010010110000000000000000;
		112: Instruction <= 32'b00100001011010110000100000000000;
		113: Instruction <= 32'b10101110001010110000000000010100;
		114: Instruction <= 32'b00000000000000000000000000000000;
		115: Instruction <= 32'b00000000000000000000000000000000;
		116: Instruction <= 32'b00000000000000000000000000000000;
		117: Instruction <= 32'b00000000000000000000000000000000;
		118: Instruction <= 32'b00111100000010010000000000000000;
		119: Instruction <= 32'b10101110001010010000000000010100;
		120: Instruction <= 32'b00111100000010100000000000000000;
		121: Instruction <= 32'b00100001010010100000000000000011;
		122: Instruction <= 32'b10101110001010100000000000001000;
		123: Instruction <= 32'b10001111101010110000000000001000;
		124: Instruction <= 32'b10001111101010100000000000000100;
		125: Instruction <= 32'b10001111101010010000000000000000;
		126: Instruction <= 32'b00100011101111010000000000001100;
		127: Instruction <= 32'b00000011010000000000000000001000;
		128: Instruction <= 32'b00000011010000000000000000001000;

		default: Instruction <= 32'h08001000;	// 
		
		endcase
		
endmodule
