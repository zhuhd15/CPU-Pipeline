module PC_Adder(PC,PCplus4);
	input PC;
	output  PCplus4;
	endmodule